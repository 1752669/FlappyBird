`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/05/23 23:24:04
// Design Name: 
// Module Name: inst
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module inst(
input [31:0] instructionCode, // 指令
    output reg [53:0] decodedData
    );
    always @(*) begin
    casex ({instructionCode[31:26], instructionCode[5:0]})
    12'b000000100000: decodedData = 54'b000000000000000000000000000000000000000000000000000001; // add
    12'b000000100001: decodedData = 54'b000000000000000000000000000000000000000000000000000010; // addu
    12'b000000100010: decodedData = 54'b000000000000000000000000000000000000000000000000000100; // sub
    12'b000000100011: decodedData = 54'b000000000000000000000000000000000000000000000000001000; // subu
    12'b000000100100: decodedData = 54'b000000000000000000000000000000000000000000000000010000; // and
    12'b000000100101: decodedData = 54'b000000000000000000000000000000000000000000000000100000; // or
    12'b000000100110: decodedData = 54'b000000000000000000000000000000000000000000000001000000; // xor
    12'b000000100111: decodedData = 54'b000000000000000000000000000000000000000000000010000000; // nor
    12'b000000101010: decodedData = 54'b000000000000000000000000000000000000000000000100000000; // slt
    12'b000000101011: decodedData = 54'b000000000000000000000000000000000000000000001000000000; // sltu
    12'b000000000000: decodedData = 54'b000000000000000000000000000000000000000000010000000000; // sll
    12'b000000000010: decodedData = 54'b000000000000000000000000000000000000000000100000000000; // srl
    12'b000000000011: decodedData = 54'b000000000000000000000000000000000000000001000000000000; // sra
    12'b000000000100: decodedData = 54'b000000000000000000000000000000000000000010000000000000; // sllv
    12'b000000000110: decodedData = 54'b000000000000000000000000000000000000000100000000000000; // srlv
    12'b000000000111: decodedData = 54'b000000000000000000000000000000000000001000000000000000; // srav
    12'b000000001000: decodedData = 54'b000000000000000000000000000000000000010000000000000000; // jr
    12'b001000xxxxxx: decodedData = 54'b000000000000000000000000000000000000100000000000000000; // addi
    12'b001001xxxxxx: decodedData = 54'b000000000000000000000000000000000001000000000000000000; // addiu
    12'b001100xxxxxx: decodedData = 54'b000000000000000000000000000000000010000000000000000000; // andi
    12'b001101xxxxxx: decodedData = 54'b000000000000000000000000000000000100000000000000000000; // ori
    12'b001110xxxxxx: decodedData = 54'b000000000000000000000000000000001000000000000000000000; // xori
    12'b100011xxxxxx: decodedData = 54'b000000000000000000000000000000010000000000000000000000; // lw
    12'b101011xxxxxx: decodedData = 54'b000000000000000000000000000000100000000000000000000000; // sw
    12'b000100xxxxxx: decodedData = 54'b000000000000000000000000000001000000000000000000000000; // beq
    12'b000101xxxxxx: decodedData = 54'b000000000000000000000000000010000000000000000000000000; // bne
    12'b001010xxxxxx: decodedData = 54'b000000000000000000000000000100000000000000000000000000; // slti
    12'b011100xxxxxx:
        if (instructionCode[5:0] == 6'b000010)
            decodedData = 54'b000000100000000000000000000000000000000000000000000000; // mul
        else
            decodedData = 54'b000000000000000000000010000000000000000000000000000000; // clz
    12'b001011xxxxxx: decodedData = 54'b000000000000000000000000001000000000000000000000000000; // sltiu
    12'b001111xxxxxx: begin
        if (instructionCode[25:21] == 5'b0)
            decodedData = 54'b000000000000000000000000010000000000000000000000000000; // lui
        else
            decodedData = 54'bz;
    end
    12'b000010xxxxxx: decodedData = 54'b000000000000000000000000100000000000000000000000000000; // j
    12'b000011xxxxxx: decodedData = 54'b000000000000000000000001000000000000000000000000000000; // jal
    12'b000000011011: decodedData = 54'b000000000000000000000100000000000000000000000000000000; // divu
    12'b010000011000: decodedData = 54'b000000000000000000001000000000000000000000000000000000; // eret
    12'b000000001001: decodedData = 54'b000000000000000000010000000000000000000000000000000000; // jalr
    12'b100000xxxxxx: decodedData = 54'b000000000000000000100000000000000000000000000000000000; // lb
    12'b100100xxxxxx: decodedData = 54'b000000000000000001000000000000000000000000000000000000; // lbu
    12'b100101xxxxxx: decodedData = 54'b000000000000000010000000000000000000000000000000000000; // lhu
    12'b101000xxxxxx: decodedData = 54'b000000000000000100000000000000000000000000000000000000; // sb
    12'b101001xxxxxx: decodedData = 54'b000000000000001000000000000000000000000000000000000000; // sh
    12'b100001xxxxxx: decodedData = 54'b000000000000010000000000000000000000000000000000000000; // lh
    12'b010000000000: 
    begin
        if (instructionCode[25:21] == 5'b00000)
            decodedData = 54'b000000000000100000000000000000000000000000000000000000; // mfc0
        else
            decodedData = 54'b000000000100000000000000000000000000000000000000000000; // mtc0
            end
    12'b000000010000: decodedData = 54'b000000000001000000000000000000000000000000000000000000; // mfh1
    12'b000000010010: decodedData = 54'b000000000010000000000000000000000000000000000000000000; // mflo
    12'b010000000000: decodedData = 54'b000000000100000000000000000000000000000000000000000000; // mtc0
    12'b000000010001: decodedData = 54'b000000001000000000000000000000000000000000000000000000; // mth1
    12'b000000010011: decodedData = 54'b000000010000000000000000000000000000000000000000000000; // mtlo
    12'b000000011001: decodedData = 54'b000001000000000000000000000000000000000000000000000000; // multu
    12'b000000001100: decodedData = 54'b000010000000000000000000000000000000000000000000000000; // syscall
    12'b000000110100: decodedData = 54'b000100000000000000000000000000000000000000000000000000; // teq
    12'b000001xxxxxx: decodedData = 54'b001000000000000000000000000000000000000000000000000000; // bgez
    12'b000000001101: decodedData = 54'b010000000000000000000000000000000000000000000000000000; // break
    12'b000000011010: decodedData = 54'b100000000000000000000000000000000000000000000000000000; // div

    default: decodedData = 54'bz;
    endcase
end

endmodule
